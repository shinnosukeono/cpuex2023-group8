module address_buffer #(
    parameter EVAL_DELAY = 2
) (
    input clk, rst,
        
);
    
endmodule