`ifndef _const_h
`define _const_h
localparam AXI_ADDRW = 4;
localparam AXI_DATAW = 32;
localparam DATAW = 32;
localparam UART_ADDR = 0;
localparam DATA_MEM_ADDR = 0;
localparam INST_MEM_ADDR = 0;
localparam INST_MEM_ADDRW = 32;
localparam CACHE_LINEW = 32;
localparam CACHE_ADDRW = 32;
`endif