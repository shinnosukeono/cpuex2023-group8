`timescale 1ps/1ps

module TEST(); //ここを名前に

reg[31:0] a;
reg[31:0] b;
wire[31:0] c;
reg[31:0] i;
integer j=3;
logic clk;
logic rst;

fsub_pipe and_instance(clk,rst,a, b, c); //オブジェクト指向感

initial begin

        a = 32'h00000000; b = 32'h00000000;
        #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0;

        for (i = 0; i < 100000; i += 1) begin
                #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0;

                #2 $display("%b %b %b", a, b, c);
                #2 a = $random(j) % 32'hFFFFFFFF;
                #2 b = $random(j) % 32'hFFFFFFFF;
        end
        #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0;

        #2 $display("%b %b %b", a, b, c);
        #2 a = 32'hFFFFFFFF; b = 32'hFFFFFFFF;
        #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0; #3 clk = 1'b1; #3 clk = 1'b0;

        #2 $display("%b %b %b", a, b, c);

        #10 $finish;
end

endmodule