module instr_gen (
    input wire clk,
    input wire [31:0] counter,
    output reg addr_sel,
    output wire we,
    output reg [31:0] addr,
    output wire [31:0] dout
);
    localparam LEN = 'd128;
    logic [31:0] instr_array [0:LEN-1];
    assign instr_array = {
        // int fib
        // 32'hfe010113,
        // 32'h00112e23,
        // 32'h00812c23,
        // 32'h02010413,
        // 32'hfe042623,
        // 32'hfe042423,
        // 32'h00100793,
        // 32'hfef42223,
        // 32'h0300006f,
        // 32'hfe442703,
        // 32'hfe842783,
        // 32'h00f707b3,
        // 32'hfef42023,
        // 32'hfe442783,
        // 32'hfef42423,
        // 32'hfe042783,
        // 32'hfef42223,
        // 32'hfec42783,
        // 32'h00178793,
        // 32'hfef42623,
        // 32'hfec42703,
        // 32'h00900793,
        // 32'hfce7d6e3,
        // 32'h00000793,
        // 32'h00078513,
        // 32'h01c12083,
        // 32'h01812403,
        // 32'h02010113,
        // 32'h000fd073

        // floating fib
        // 32'h3f8007b7,
        // 32'h06f02c23,
        // 32'hfe010113,
        // 32'h00112e23,
        // 32'h00812c23,
        // 32'h02010413,
        // 32'hfe042623,
        // 32'hfe042423,
        // 32'h000007b7,
        // 32'h0807a787,
        // 32'hfef42227,
        // 32'h0300006f,
        // 32'hfe442707,
        // 32'hfe842787,
        // 32'h00f777d3,
        // 32'hfef42027,
        // 32'hfe442787,
        // 32'hfef42427,
        // 32'hfe042787,
        // 32'hfef42227,
        // 32'hfec42783,
        // 32'h00178793,
        // 32'hfef42623,
        // 32'hfec42703,
        // 32'h00900793,
        // 32'hfce7d6e3,
        // 32'h00000793,
        // 32'h00078513,
        // 32'h01c12083,
        // 32'h01812403,
        // 32'h02010113,
        // 32'h000fd073

        // int fib recursive
        // 32'hfe010113,
        // 32'h00112e23,
        // 32'h00812c23,
        // 32'h02010413,
        // 32'h00a00513,
        // 32'h028000ef,
        // 32'hfea42623,
        // 32'hfec42583,
        // 32'h00058013,
        // 32'h00000793,
        // 32'h00078513,
        // 32'h01c12083,
        // 32'h01812403,
        // 32'h02010113,
        // 32'h000fd073,
        // 32'hfe010113,
        // 32'h00112e23,
        // 32'h00812c23,
        // 32'h02010413,
        // 32'hfea42623,
        // 32'hfec42783,
        // 32'h00179793,
        // 32'h00078513,
        // 32'h01c12083,
        // 32'h01812403,
        // 32'h02010113,
        // 32'h00008067
32'hfe010113,
32'h00112e23,
32'h00812c23,
32'h02010413,
32'h000107b7,
32'h0007a787,
32'hfef42627,
32'h000107b7,
32'h0047a787,
32'h20f785d3,
32'hfec42507,
32'h028000ef,
32'hfea42427,
32'hfe842507,
32'h0c4000ef,
32'h00000793,
32'h00078513,
32'h01c12083,
32'h01812403,
32'h02010113,
32'h000fd073,
32'hfd010113,
32'h02112623,
32'h02812423,
32'h03010413,
32'hfca42e27,
32'hfcb42c27,
32'hfdc42707,
32'h000107b7,
32'h0007a787,
32'h18f777d3,
32'hfef42627,
32'h0280006f,
32'hfdc42707,
32'hfec42787,
32'h18f77753,
32'hfec42787,
32'h00f77753,
32'h000107b7,
32'h0087a787,
32'h10f777d3,
32'hfef42627,
32'hfec42787,
32'h10f7f753,
32'hfdc42787,
32'h08f777d3,
32'hfd842707,
32'ha0f717d3,
32'hfc0792e3,
32'hfec42787,
32'h10f7f753,
32'hfdc42787,
32'h08f77753,
32'hfd842787,
32'h20f797d3,
32'ha0f717d3,
32'hfa0792e3,
32'hfec42787,
32'h20f78553,
32'h02c12083,
32'h02812403,
32'h03010113,
32'h00008067,
32'hfd010113,
32'h02112623,
32'h02812423,
32'h03010413,
32'hfca42e27,
32'hfdc40793,
32'hfef42423,
32'hfe842783,
32'h0007a783,
32'hfef42223,
32'h01f00793,
32'hfef42623,
32'h0380006f,
32'hfec42783,
32'hfe442703,
32'h00f757b3,
32'h0017f793,
32'h00078663,
32'h03100793,
32'h0080006f,
32'h03000793,
32'h00078513,
32'h034000ef,
32'hfec42783,
32'hfff78793,
32'hfef42623,
32'hfec42783,
32'hfc07d4e3,
32'h00a00513,
32'h018000ef,
32'h00000013,
32'h02c12083,
32'h02812403,
32'h03010113,
32'h00008067,
32'h00050011,
32'h00008067
    };

    always @(posedge clk) begin
        addr_sel <= we;
    end

    assign we = (counter <= 32'h80) ? 1'b1 : 1'b0;

    always @(posedge clk) begin
        if (counter == 32'h80) begin
            addr <= 32'b0;
        end
        else if (counter < 32'h80) begin
            addr <= (counter >> 2) << 2;
        end
    end

    assign dout = ((addr>>2) < 'd128) ? instr_array[(addr >> 2)] : 32'b0;
endmodule