`ifndef _io_params_vh_
`define _io_params_vh_
// parameter _CLK_PER_HALF_BIT = 108;  // 50,000,000 (Hz) / (230400 (baudrate) * 2)
parameter _CLK_PER_HALF_BIT = 174;  // 80,200,000 (MHz) / (230,400 (baudrate) * 2)
// parameter _CLK_PER_HALF_BIT = 2607;  // 50,000,000 (Hz) / (9600 (baudrate) * 2)
`endif