`ifndef _io_params_vh_
`define _io_params_vh_
parameter _CLK_PER_HALF_BIT = 217;  // 50,000,000 (MHz) / (115,200 (baudrate) * 2)
`endif