module test_wrapper (
    input wire clk
);
    test i_test (
        .clk(clk)
    );
endmodule